library ieee;
use ieee.std_logic_1164.all;

library work;
use work.std_logic_vector_to_string_package.all;

entity alu_tb is
--  A testbench has no ports.
end alu_tb;

architecture behaviour of alu_tb is
	--  Declaration of the component that will be instantiated.
	component alu
		port (
			x  : in std_logic_vector(0 to 15);
			y  : in std_logic_vector(0 to 15);
			zx : in std_logic;                  
			nx : in std_logic;
			zy : in std_logic;
			ny : in std_logic;
			f  : in std_logic;
			no : in std_logic;
	
			out0 : out std_logic_vector(0 to 15);
			zr : out std_logic;
			ng : out std_logic
		);
  	end component;

	--  Specifies which entity is bound with the component.
	for alu_0: alu use entity work.alu;
	signal x, y, out0 : std_logic_vector(0 to 15);
	signal zx, nx, zy, ny, f, no, zr, ng : std_logic;

begin
	--  Component instantiation.
	alu_0: alu port map (
		x => x,
		y => y,
		zx => zx,                  
		nx => nx,
		zy => zy,
		ny => ny,
		f  => f,
		no => no,

		out0 => out0,
		zr => zr,
		ng => ng
	);

	--  This process does the real job.
	process
		type pattern_type is record
			--  The inputs.
			x, y : std_logic_vector(0 to 15);
			zx, nx, zy, ny, f, no : std_logic;
			--  The expected outputs.
			out0 : std_logic_vector(0 to 15);
			zr, ng : std_logic;			
		end record;

		--  The patterns to apply.
		type pattern_array is array (natural range <>) of pattern_type;
		constant patterns : pattern_array :=
		(			
			("0000000000000000", "1111111111111111", '1', '0', '1', '0', '1', '0', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '1', '1', '1', '1', "1000000000000000", '0', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '1', '0', '1', '0', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '0', '1', '1', '0', '0', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '0', '0', '0', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '0', '1', '1', '0', '1', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '0', '0', '1', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '0', '0', '1', '1', '1', '1', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '0', '1', '1', "1000000000000000", '0', '0'),
			("0000000000000000", "1111111111111111", '0', '1', '1', '1', '1', '1', "1000000000000000", '0', '0'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '1', '1', '1', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '0', '0', '1', '1', '1', '0', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '1', '1', '0', '0', '1', '0', "0111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '0', '0', '0', '1', '0', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '1', '0', '0', '1', '1', "1000000000000000", '0', '0'),
			("0000000000000000", "1111111111111111", '0', '0', '0', '1', '1', '1', "1111111111111111", '0', '1'),
			("0000000000000000", "1111111111111111", '0', '0', '0', '0', '0', '0', "0000000000000000", '1', '0'),
			("0000000000000000", "1111111111111111", '0', '1', '0', '1', '0', '1', "1111111111111111", '0', '1'),
			("1000100000000000", "1100000000000000", '1', '0', '1', '0', '1', '0', "0000000000000000", '1', '0'),
			("1000100000000000", "1100000000000000", '1', '1', '1', '1', '1', '1', "1000000000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '1', '1', '1', '0', '1', '0', "1111111111111111", '0', '1'),
			("1000100000000000", "1100000000000000", '0', '0', '1', '1', '0', '0', "1000100000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '1', '1', '0', '0', '0', '0', "1100000000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '0', '0', '1', '1', '0', '1', "0111011111111111", '0', '1'),
			("1000100000000000", "1100000000000000", '1', '1', '0', '0', '0', '1', "0011111111111111", '0', '1'),
			("1000100000000000", "1100000000000000", '0', '0', '1', '1', '1', '1', "1111011111111111", '0', '1'),
			("1000100000000000", "1100000000000000", '1', '1', '0', '0', '1', '1', "1011111111111111", '0', '1'),
			("1000100000000000", "1100000000000000", '0', '1', '1', '1', '1', '1', "0100100000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '1', '1', '0', '1', '1', '1', "0010000000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '0', '0', '1', '1', '1', '0', "0000100000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '1', '1', '0', '0', '1', '0', "0100000000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '0', '0', '0', '0', '1', '0', "0010100000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '0', '1', '0', '0', '1', '1', "0111000000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '0', '0', '0', '1', '1', '1', "0100111111111111", '0', '1'),
			("1000100000000000", "1100000000000000", '0', '0', '0', '0', '0', '0', "1000000000000000", '0', '0'),
			("1000100000000000", "1100000000000000", '0', '1', '0', '1', '0', '1', "1100100000000000", '0', '0')			
		);
	begin
		--  Check each pattern.
		for i in patterns'range loop
			--  Set the inputs.
			x <= patterns(i).x;
			y <= patterns(i).y;
			zx <= patterns(i).zx;
			nx <= patterns(i).nx;
			zy <= patterns(i).zy;
			ny <= patterns(i).ny;
			f <= patterns(i).f;
			no <= patterns(i).no;			
			--  Wait for the results.
			wait for 1 ns;
			--  Check the outputs.
			assert out0 = patterns(i).out0
			report "bad value for i = " & integer'image(i)
					& " out0 " & to_string(out0) & " instead of " & to_string(patterns(i).out0)
			severity error;
			
			assert zr = patterns(i).zr
			report "bad value for i = " & integer'image(i)
					& " zr " & std_logic'image(zr) & " instead of " & std_logic'image(patterns(i).zr)
			severity error;
			
			assert ng = patterns(i).ng						
			report "bad value for i = " & integer'image(i)
					& " ng " & std_logic'image(ng) & " instead of " & std_logic'image(patterns(i).ng)									
			severity error;
		end loop;

		assert false report "end of test" severity note;
		--  Wait forever; this will finish the simulation.
		wait;
	end process;

end behaviour;
