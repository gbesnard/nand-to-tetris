library ieee;
use ieee.std_logic_1164.all;

entity mux8way16_gate_tb is
--  A testbench has no ports.
end mux8way16_gate_tb;

architecture behaviour of mux8way16_gate_tb is
	--  Declaration of the component that will be instantiated.
	component mux8way16_gate
		port (
			in0 : in std_logic_vector(0 to 15);
			in1 : in std_logic_vector(0 to 15);
			in2 : in std_logic_vector(0 to 15);
			in3 : in std_logic_vector(0 to 15);
			in4 : in std_logic_vector(0 to 15);
			in5 : in std_logic_vector(0 to 15);
			in6 :  std_logic_vector(0 to 15);
			in7 :  std_logic_vector(0 to 15); 
			sel0 : in std_logic_vector(0 to 2); 
			out0 : out std_logic_vector(0 to 15)

		);
  	end component;

	--  Specifies which entity is bound with the component.
	for mux8way16_gate_0: mux8way16_gate use entity work.mux8way16_gate;
	signal in0, in1, in2, in3, in4, in5, in6, in7, out0 : std_logic_vector(0 to 15);
	signal sel0 : std_logic_vector(0 to 2);

begin
	--  Component instantiation.
	mux8way16_gate_0: mux8way16_gate port map (
		in0 => in0, 
		in1 => in1, 
		in2 => in2, 
		in3 => in3, 
		in4 => in4, 
		in5 => in5, 
		in6 => in6, 
		in7 => in7, 
		sel0 => sel0, 
		out0 => out0
	);

	--  This process does the real job.
	process
		type pattern_type is record
			--  The inputs of the mux8way16_gate.
			in0 : std_logic_vector(0 to 15);
			in1 : std_logic_vector(0 to 15);
			in2 : std_logic_vector(0 to 15);
			in3 : std_logic_vector(0 to 15);
			in4 : std_logic_vector(0 to 15);
            in5 : std_logic_vector(0 to 15);
            in6 : std_logic_vector(0 to 15);
            in7 : std_logic_vector(0 to 15);
            sel0 : std_logic_vector(0 to 2);
			--  The expected outputs of the adder.
			out0 : std_logic_vector(0 to 15);
		end record;

		--  The patterns to apply.
		type pattern_array is array (natural range <>) of pattern_type;
		constant patterns : pattern_array :=
		(
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "000", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "001", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "010", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "011", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "100", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "101", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "110", "0000000000000000"),
			("0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "111", "0000000000000000"),

			("0001001000110100", "0010001101000101", "0011010001010110", "0100010101100111", "0101011001111000", "0110011110001001", "0111100010011010", "1000100110101011", "000", "0001001000110100"),
			("0001001000110100", "0010001101000101", "0011010001010110", "0100010101100111", "0101011001111000", "0110011110001001", "0111100010011010", "1000100110101011", "001", "0101011001111000"),
			("0001001000110100", "0010001101000101", "0011010001010110", "0100010101100111", "0101011001111000", "0110011110001001", "0111100010011010", "1000100110101011", "010", "0011010001010110"),
			("0001001000110100", "0010001101000101", "0011010001010110", "0100010101100111", "0101011001111000", "0110011110001001", "0111100010011010", "1000100110101011", "011", "0111100010011010"),
			("0001001000110100", "0010001101000101", "0011010001010110", "0100010101100111", "0101011001111000", "0110011110001001", "0111100010011010", "1000100110101011", "100", "0010001101000101"),
			("0001001000110100", "0010001101000101", "0011010001010110", "0100010101100111", "0101011001111000", "0110011110001001", "0111100010011010", "1000100110101011", "101", "0110011110001001"),
			("0001001000110100", "0010001101000101", "0011010001010110", "0100010101100111", "0101011001111000", "0110011110001001", "0111100010011010", "1000100110101011", "110", "0100010101100111"),
			("0001001000110100", "0010001101000101", "0011010001010110", "0100010101100111", "0101011001111000", "0110011110001001", "0111100010011010", "1000100110101011", "111", "1000100110101011")
		);

	begin
		--  Check each pattern.
		for i in patterns'range loop

			--  Set the inputs.
			in0 <= patterns(i).in0;
			in1 <= patterns(i).in1;
			in2 <= patterns(i).in2;
			in3 <= patterns(i).in3;
			in4 <= patterns(i).in4;
			in5 <= patterns(i).in5;
			in6 <= patterns(i).in6;
			in7 <= patterns(i).in7;
			sel0 <= patterns(i).sel0;
			--  Wait for the results.
			wait for 1 ns;
			--  Check the outputs.
			assert out0 = patterns(i).out0
			report "bad value" severity error;
		end loop;

		assert false report "end of test" severity note;
		--  Wait forever; this will finish the simulation.
		wait;
	end process;

end behaviour;
